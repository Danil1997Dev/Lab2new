// niosII_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module niosII_tb (
	);

	wire    niosii_inst_clk_bfm_clk_clk;       // niosII_inst_clk_bfm:clk -> [niosII_inst:clk_clk, niosII_inst_reset_bfm:clk]
	wire    niosii_inst_reset_bfm_reset_reset; // niosII_inst_reset_bfm:reset -> niosII_inst:reset_reset_n
	reg train;
	wire red, yellow, green;

	niosII niosii_inst (
		.clk_clk           (niosii_inst_clk_bfm_clk_clk),       //        clk.clk
		.reset_reset_n     (niosii_inst_reset_bfm_reset_reset), //      reset.reset_n
		.sem_export_train  (train),                                  // sem_export.train
		.sem_export_red    (red),                                  //           .red
		.sem_export_yellow (yellow),                                  //           .yellow
		.sem_export_green  (green)                                   //           .green
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) niosii_inst_clk_bfm (
		.clk (niosii_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) niosii_inst_reset_bfm (
		.reset (niosii_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (niosii_inst_clk_bfm_clk_clk)        //   clk.clk
	);
	
	initial
	begin
$monitor("divider = %b", niosii_inst.sem.divider) ;  
		train = 0;
		wait (niosii_inst_reset_bfm_reset_reset);
		forever
		begin
			repeat(16000)@(posedge niosii_inst_clk_bfm_clk_clk);
			train = 1;
			repeat(10)@(posedge niosii_inst_clk_bfm_clk_clk);
			train = 0;
		end
	end

endmodule
